module Four(out);

	output reg [31:0] out;
	
	always begin
		out = 4;
	end

endmodule 